// Copyright (C) 1991-2004 Altera Corporation
// Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
// support information,  device programming or simulation file,  and any other
// associated  documentation or information  provided by  Altera  or a partner
// under  Altera's   Megafunction   Partnership   Program  may  be  used  only
// to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
// other  use  of such  megafunction  design,  netlist,  support  information,
// device programming or simulation file,  or any other  related documentation
// or information  is prohibited  for  any  other purpose,  including, but not
// limited to  modification,  reverse engineering,  de-compiling, or use  with
// any other  silicon devices,  unless such use is  explicitly  licensed under
// a separate agreement with  Altera  or a megafunction partner.  Title to the
// intellectual property,  including patents,  copyrights,  trademarks,  trade
// secrets,  or maskworks,  embodied in any such megafunction design, netlist,
// support  information,  device programming or simulation file,  or any other
// related documentation or information provided by  Altera  or a megafunction
// partner, remains with Altera, the megafunction partner, or their respective
// licensors. No other licenses, including any licenses needed under any third
// party's intellectual property, are provided herein.

module TOP(
	In_Wen,
	In_Wclk,
	In_Rclk,
	In_Raddr,
	In_Waddr,
	In_Wdata,
	Out_Rdata
);

input	In_Wen;
input	In_Wclk;
input	In_Rclk;
input	[4:0] In_Raddr;
input	[4:0] In_Waddr;
input	[7:0] In_Wdata;
output	[7:0] Out_Rdata;






DualPortRAM	b2v_inst(.wren(In_Wen),.wrclock(In_Wclk),.rdclock(In_Rclk),.data(In_Wdata),.rdaddress(In_Raddr),.wraddress(In_Waddr),.q(Out_Rdata));


endmodule
